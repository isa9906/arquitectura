library IEEE;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity codificando is
	port
	(
		-- Input ports
		x1	: in  std_logic;
		x2	: in  std_logic;
		x3	: in  std_logic;
		x4	: in  std_logic;
		x5	: in  std_logic;
		x6	: in  std_logic;
		x7	: in  std_logic;
		x8	: in  std_logic;
		x9	: in  std_logic;
		x0	: in  std_logic;
		

		

		-- Output ports
		a	: out  std_logic;
		b	: out  std_logic;
		c	: out  std_logic;
		d	: out  std_logic
	);
end codificando;

architecture comportamiento of codificando is

	

begin

	a<= (x8 or x9);
	b<= (x4 or x5 or x6 or x7);
	c<= (x2 or x3 or x6 or x7);
	d<= (x1 or x3 or x5 or x7 or x9);
	-- esta es extraida de la tabla de verdad. 

end comportamiento;

